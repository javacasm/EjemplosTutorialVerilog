//------------------------------------------------------------------
//-- Verilog template
//-- Top entity
//-- Board: icezum
//------------------------------------------------------------------
`default_nettype none

//-- Fichero setbit.v
module setbit(output A);
wire A;

assign A = 1;

endmodule
